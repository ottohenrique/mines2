[[o:	Cell:@valueI"1:EF:@state:playedo; ;I"x;T;:closedo; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	[o; ;I"1;F;;
o; ;I"1;F;;
o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I"1;F;;	[o; ;I" ;T;;
o; ;I"1;F;;
o; ;I"1;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"x;T;:flaggedo; ;I"1;F;;
[o; ;I" ;T;;
o; ;I"1;F;;
o; ;I"x;T;;
o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I"1;F;;	[o; ;I" ;T;;
o; ;I"1;F;;
o; ;I"2;F;;
o; ;I"2;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"2;F;;	o; ;I"2;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"x;T;;
o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	[o; ;I" ;T;;
o; ;I" ;T;;
o; ;I"1;F;;
o; ;I"x;T;;
o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"2;F;;	o; ;I"x;T;;
o; ;I"x;T;;
o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	[o; ;I"1;F;;
o; ;I"1;F;;
o; ;I"2;F;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"2;F;;	o; ;I"x;T;;
o; ;I"3;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	[o; ;I"1;F;;
o; ;I"x;T;;o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"x;T;;
o; ;I"2;F;;	o; ;I"1;F;;	o; ;I" ;T;;	[o; ;I"1;F;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"2;F;;	o; ;I"2;F;;	o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"1;F;;	o; ;I"3;F;;	o; ;I"3;F;;
o; ;I"x;T;;
o; ;I"1;F;;	o; ;I" ;T;;	[o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"x;T;;
o; ;I"x;T;;
o; ;I"1;F;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I" ;T;;	o; ;I"1;F;;	o; ;I"x;T;;
o; ;I"2;F;;
o; ;I"x;T;;
o; ;I"2;F;;
o; ;I"1;F;;	o; ;I" ;T;;	